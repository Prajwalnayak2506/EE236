Shunt Clipper DC analysis
r1 1 2 1k
*Specifying a default diode p n
d1 2 3 di
.model di D()
*Independent DC source of 2V
vdc 0 3 dc 2
*Independent DC source whose voltage is to be varied
vin 1 0 sin (0 5v 1k 0 0)
.tran 0.01m 6m
.control
run
plot v(1) v(2)
.endc
