All in one figures
*including the txts
.include rn142.txt

*Diode
r0  gnd 2 500
c0  1 2 100n
v_1 20 2 dc 0
d0  3 20 DRN142S
r1  6 3 500
c1  3 4 100n
r2  4 40 50
v_2 40 gnd dc 0

vbias gnd 6 dc 0
vin gnd 1 sin (0 6V 1Meg 0 0)
*DC Analysis on source vin, to vary from 0 to +5V
.tran 0.1n 3u
.control
* Define values of vbias and corresponding filenames
let bias_values = [-5, 0, 1, 3, 5]
let filenames = ["voltages_bias_-5V.ps", "voltages_bias_0V.ps", "voltages_bias_1V.ps", "voltages_bias_3V.ps", "voltages_bias_5V.ps"]
let current_filenames = ["currents_bias_-5V.ps", "currents_bias_0V.ps", "currents_bias_1V.ps", "currents_bias_3V.ps", "currents_bias_5V.ps"]

* Iterate over bias values
let i = 0
foreach val bias_values
    alter vbias dc val
    run
    * Use filenames array to save plots
    plot v(1) v(4)
    set hcopydevtype=postscript
    hardcopy C:\Users\Public\filenames[i] v(1) v(4)
    plot I(v_1) I(v_2)
    hardcopy C:\Users\Public\current_filenames[i] I(v_1) I(v_2)
    let i = i + 1
end
.endc
.end
