 Diode I-V characteristics
*Including the predefined op-amp subcircuit file
.include white_5mm.txt
*Connections as mentioned in subcircuit file
d1 1 2 WHITE
r1 2 0 100
v1 1 0 12
.control
run
dc V1 0.0001 5 0.0001
plot -i(V1)
plot ln(-i(V1))
.endc
.end

