5 in one
.include white_5mm.txt
.include red_5mm.txt
.include blue_5mm.txt
.include green_5mm.txt
.include PN_1N4007.txt

r1 2 3 100
v1 3 0 dc 0

r2 6 66 100
v2 66 0 dc 0

r3 7 77 100
v3 77 0 dc 0

r4 8 88 100
v4 88 0 dc 0

r5 9 99 100
v5 99 0 dc 0

d1 1 2 BLUE
d2 1 6 WHITE
d3 1 7 GREEN
d4 1 8 RED
d5 1 9 1N4007

vin 1 0 dc 0
.dc vin 0.1 5 0.01
.control
run
let vd = v(1) - v(2)
plot ln(i(v1)) vs vd  ln(i(v2)) vs v(1)-v(6)  ln(i(v3)) vs v(1)-v(7)  ln(i(v4)) vs v(1)-v(8)  ln(i(v5)) vs v(1)-v(9)
plot i(v1) vs vd  i(v2) vs v(1)-v(6)  i(v3) vs v(1)-v(7)  i(v4) vs v(1)-v(8)  i(v5) vs v(1)-v(9)


 .endc
 .end